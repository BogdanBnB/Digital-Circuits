`timescale 1ns / 1ps

module Half_adder(
        input in0,
        input in1
    );
assign {cout,out0}=in0+in1;
endmodule
