`timescale 1ns / 1ps
module sumator(
        input in0,
        input in1
    );

assign out=in0+in1;
endmodule
